module data_sw(
							clk,
							res,
							data_in,
							data_in_comp,
							sw,
							data_out
							);
input 					clk,res;//ʱ�Ӻ͸�λ��
input[7:0]				data_in,data_in_comp;//����ԭ��Ͳ������룻
input					sw;//ԭ�벹���л���
output[7:0]			data_out;//���������

reg[7:0]				data_out;

always@(posedge clk or negedge res) 
if(!res) begin
	data_out<=0;
end
else begin
	data_out<=sw?data_in_comp:data_in;//ԭ�벹���л���
end
endmodule
