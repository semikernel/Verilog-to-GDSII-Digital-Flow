module data_pro(
							clk,
							res,
							data_in_a,
							data_in_b,
							en_data_in,
							data_out,
							data_out_comp,
							en_data_out
							);
input 					clk,res;//ʱ�Ӻ͸�λ��
input[3:0]				data_in_a,data_in_b;//�������룻
input					en_data_in;//��������ʹ�ܣ�
output[7:0]			data_out,data_out_comp;//����ԭ��Ͳ��������
input					en_data_out;//�������ʹ�ܣ�

reg[3:0]				buf_a,buf_b;//��������Ĵ�����
reg[3:0]				buf_a_dealy,buf_b_dealy;//��ʱһ�ļĴ�����
reg[7:0]				data_out;

//����ת����
assign					data_out_comp=data_out[7]?{data_out[7],~data_out[6:0]+1}:data_out;

always@(posedge clk or negedge res) 
if(!res) begin
	buf_a<=0;buf_b<=0;
	buf_a_dealy<=0;buf_b_dealy<=0;
	data_out<=0;
end
else begin
	//�������벢��1��
	if(en_data_in) begin
		buf_a<=data_in_a+1;
		buf_b<=data_in_b+1;
	end
	//��ʱһ�ģ�
	buf_a_dealy<=buf_a;
	buf_b_dealy<=buf_b;
	//�˷����㣻
	if(en_data_out) begin
		data_out<=buf_a_dealy*buf_b_dealy;
	end	
end
endmodule



